library verilog;
use verilog.vl_types.all;
entity RIPPLECOUNTER_vlg_vec_tst is
end RIPPLECOUNTER_vlg_vec_tst;
